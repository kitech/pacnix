module main

fn test_1() {}

fn test_2() {

	assert false
}